//sample6.v 1







//sample.v 1


module sample ;
    wire out;
    assign out=1;

endmodule


//sample6.v 8


module sample2 ;
    wire out;
    assign out=1;

endmodule


