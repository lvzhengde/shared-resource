`define X 1

module sample ;
    wire out ;
    assign out=`X;

endmodule

