//sample2.v 1


module sample ;
    wire out;
    assign out=1;

endmodule


