module sample1 ;
    parameter XXX=1;
    wire out;
    assign out=XXX;
endmodule



