
`include "sample.v"
module sample2 ;
    wire out;
    assign out=1;

endmodule

