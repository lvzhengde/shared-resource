//sample9.v 1


























module sample2 ;
    wire out;
    assign out=1;
endmodule




