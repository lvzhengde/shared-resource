//sample7.v 1








module sample1 ;
    wire out;
    assign out=1;
endmodule













