module sample ;
    wire a;   
    wire b[1:0];
    wire[1:0] c;
    wire[1:0] d[1:0];
    wire[1:0] e[1:0],f;
    wire[1:0] g[1:0],h[1:0];
    wire[32-1:0] i[32-1:0];
    reg    j;
    input  k;
    output l;
endmodule

