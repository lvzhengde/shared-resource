`define X(n) out=n

module sample ;
    wire out;
    assign `X((1));

endmodule

