/*
    Created by Sister.
*/
module test_typedef(
    out,
    in);

    reg[1:0] proc_state_000000;
    reg[23:0] c__000001;
    reg[23:0] a__000002;
    reg[23:0] b__000002;
    reg[5:0] a__000001;
    reg[5:0] b__000001;
    reg[63:0] n;
    reg[63:0] m;
    reg[63:0] l[0:1];
    reg[63:0] k[0:1];
    reg[23:0] j;
    reg[23:0] i;
    reg[23:0] h;
    reg[5:0] g;
    reg[5:0] f;
    reg[5:0] e;
    reg[47:0] d;
    reg[23:0] c;
    reg[47:0] b;
    reg[63:0] a;
    reg[5:0] sig;
    output out;
    reg out;
    input in;

    always@( in) begin
        case(proc_state_000000)
        0 : begin
            l[1]<=170;
            l[0]<=160;
            k[1]<=150;
            k[0]<=140;
            i[23:16]<=130;
            i[15:8]<=120;
            i[7:0]<=110;
            h[23:16]<=100;
            h[15:8]<=90;
            h[7:0]<=80;
            f<=70;
            e<=60;
            d[47:40]<=50;
            c[23:16]<=40;
            c[15:8]<=30;
            b[7:0]<=20;
            a<=10;
            proc_state_000000<=1;
        end
        1 : begin
            sig<=e;
            m<=(k[0]+l[1][2:1]);
            l[1][5:3]<=190;
            k[1]<=180;
            a__000002<=h;
            b__000002<=i;
            a__000001<=e;
            b__000001<=f;
            proc_state_000000<=2;
        end
        2 : begin
            l[1][4:2]<=190;
            c__000001[23:16]<=(a__000002[23:16]+b__000002[23:16]);
            c__000001[15:8]<=(a__000002[15:8]+b__000002[15:8]);
            c__000001[7:0]<=(a__000002[7:0]+b__000002[7:0]);
            g<=(a__000001+b__000001);
            proc_state_000000<=3;
        end
        3 : begin
            n<=(k[1]+l[1]);
            m<=(k[0]+l[1][2:1]);
            j<=c__000001;
            proc_state_000000<=0;
        end
        endcase
    end

endmodule

