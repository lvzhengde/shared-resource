//sample5.v 1

//sample.v 1


module sample ;
    wire out;
    assign out=1;

endmodule


//sample5.v 2

module sample2 ;
    wire out;
    assign out=1;

endmodule


