//sample12.v 1









module sample1 ;
    wire out;
    assign out=1;
endmodule













module sample2 ;
    wire out;
    assign out=1;
endmodule



