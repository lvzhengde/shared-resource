`define X(n) n=1

module sample ;
    wire out;
    assign `X(out);

endmodule

